// display class

class display;

endclass 